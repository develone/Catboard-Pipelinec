-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity work_0CLK_83e31706 is
port(
 inputs : in work_inputs_t;
 return_output : out work_outputs_t);
end work_0CLK_83e31706;
architecture arch of work_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_efd1]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_5fac]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_a698]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_e556]
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_0b9e]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_756b]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_f197]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_2465]
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output : signed(16 downto 0);

function CONST_REF_RD_work_outputs_t_work_outputs_t_c871( ref_toks_0 : signed;
 ref_toks_1 : signed;
 ref_toks_2 : signed;
 ref_toks_3 : signed) return work_outputs_t is
 
  variable base : work_outputs_t; 
  variable return_output : work_outputs_t;
begin
      base.result(0)(0) := ref_toks_0;
      base.result(0)(1) := ref_toks_1;
      base.result(1)(0) := ref_toks_2;
      base.result(1)(1) := ref_toks_3;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right,
FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output);

-- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465 : 0 clocks latency
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right,
FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 inputs,
 -- All submodule outputs
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output,
 FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : work_outputs_t;
 variable VAR_inputs : work_inputs_t;
 variable VAR_outputs : work_outputs_t;
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_j : unsigned(31 downto 0);
 variable VAR_k : unsigned(31 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_0_0_work_h_l67_c13_9cd3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_0_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_0_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_0_1_work_h_l67_c13_9cd3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_1_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_1_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_1_0_work_h_l67_c13_9cd3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_0_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_0_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_1_1_work_h_l67_c13_9cd3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_1_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_1_work_h_l70_c17_dbc3 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output : signed(16 downto 0);
 variable VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_8985_return_output : work_outputs_t;
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_93d5_DUPLICATE_353d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_e058_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_93d5_DUPLICATE_0def_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_0b95_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_174d_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_8fac_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_93d5_DUPLICATE_3721_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_93d5_DUPLICATE_30e4_return_output : signed(7 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_1_0_work_h_l67_c13_9cd3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_1_0_work_h_l67_c13_9cd3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_0_0_work_h_l67_c13_9cd3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_outputs_result_0_0_work_h_l67_c13_9cd3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_1_1_work_h_l67_c13_9cd3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_1_1_work_h_l67_c13_9cd3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_0_1_work_h_l67_c13_9cd3 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_outputs_result_0_1_work_h_l67_c13_9cd3;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_inputs := inputs;

     -- Submodule level 0
     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d[work_h_l70_c41_93d5]_DUPLICATE_353d LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_93d5_DUPLICATE_353d_return_output := VAR_inputs.matrix0(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d[work_h_l70_c41_93d5]_DUPLICATE_0def LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_93d5_DUPLICATE_0def_return_output := VAR_inputs.matrix0(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d[work_h_l70_c41_93d5]_DUPLICATE_30e4 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_93d5_DUPLICATE_30e4_return_output := VAR_inputs.matrix0(1)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d[work_h_l70_c64_5b9c]_DUPLICATE_174d LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_174d_return_output := VAR_inputs.matrix1(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d[work_h_l70_c41_93d5]_DUPLICATE_3721 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_93d5_DUPLICATE_3721_return_output := VAR_inputs.matrix0(1)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d[work_h_l70_c64_5b9c]_DUPLICATE_e058 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_e058_return_output := VAR_inputs.matrix1(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d[work_h_l70_c64_5b9c]_DUPLICATE_8fac LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_8fac_return_output := VAR_inputs.matrix1(1)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d[work_h_l70_c64_5b9c]_DUPLICATE_0b95 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_0b95_return_output := VAR_inputs.matrix1(1)(0);

     -- Submodule level 1
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_93d5_DUPLICATE_353d_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_93d5_DUPLICATE_353d_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_93d5_DUPLICATE_0def_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_93d5_DUPLICATE_0def_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_93d5_DUPLICATE_3721_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_93d5_DUPLICATE_3721_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_93d5_DUPLICATE_30e4_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_93d5_DUPLICATE_30e4_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_e058_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_e058_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_174d_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_174d_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_0b95_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_5b9c_DUPLICATE_0b95_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_8fac_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_5b9c_DUPLICATE_8fac_return_output;
     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_7465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;

     -- Submodule level 2
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_7465_return_output;
     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_a698] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_f197] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_0b9e] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS[work_h_l70_c17_efd1] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output;

     -- Submodule level 3
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_0_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_efd1_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_1_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_a698_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_0_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0b9e_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_1_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f197_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_0_work_h_l70_c17_dbc3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_0_1_work_h_l70_c17_dbc3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_0_work_h_l70_c17_dbc3;
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left := VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_0_outputs_result_1_1_work_h_l70_c17_dbc3;
     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_756b] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_2465] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_left;
     FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output := FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_e556] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output;

     -- FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS[work_h_l70_c17_5fac] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_left;
     FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right <= VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output := FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output;

     -- Submodule level 4
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_0_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_5fac_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_1_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_e556_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_0_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_756b_return_output, 8);
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_1_work_h_l70_c17_dbc3 := resize(VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_BIN_OP_PLUS_work_h_l70_c17_2465_return_output, 8);
     -- CONST_REF_RD_work_outputs_t_work_outputs_t_c871[work_h_l74_c12_8985] LATENCY=0
     VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_8985_return_output := CONST_REF_RD_work_outputs_t_work_outputs_t_c871(
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_0_work_h_l70_c17_dbc3,
     VAR_FOR_work_h_l63_c5_1a8e_ITER_0_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_0_1_work_h_l70_c17_dbc3,
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_0_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_0_work_h_l70_c17_dbc3,
     VAR_FOR_work_h_l63_c5_1a8e_ITER_1_FOR_work_h_l65_c9_2f18_ITER_1_FOR_work_h_l68_c13_4472_ITER_1_outputs_result_1_1_work_h_l70_c17_dbc3);

     -- Submodule level 5
     VAR_return_output := VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_8985_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
