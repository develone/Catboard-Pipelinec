-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 19
entity uint32_mux16_0CLK_4e6656cf is
port(
 sel : in unsigned(3 downto 0);
 in0 : in unsigned(31 downto 0);
 in1 : in unsigned(31 downto 0);
 in2 : in unsigned(31 downto 0);
 in3 : in unsigned(31 downto 0);
 in4 : in unsigned(31 downto 0);
 in5 : in unsigned(31 downto 0);
 in6 : in unsigned(31 downto 0);
 in7 : in unsigned(31 downto 0);
 in8 : in unsigned(31 downto 0);
 in9 : in unsigned(31 downto 0);
 in10 : in unsigned(31 downto 0);
 in11 : in unsigned(31 downto 0);
 in12 : in unsigned(31 downto 0);
 in13 : in unsigned(31 downto 0);
 in14 : in unsigned(31 downto 0);
 in15 : in unsigned(31 downto 0);
 return_output : out unsigned(31 downto 0));
end uint32_mux16_0CLK_4e6656cf;
architecture arch of uint32_mux16_0CLK_4e6656cf is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- layer0_node0_MUX[bit_math_h_l18_c3_2607]
signal layer0_node0_MUX_bit_math_h_l18_c3_2607_cond : unsigned(0 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue : unsigned(31 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse : unsigned(31 downto 0);
signal layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output : unsigned(31 downto 0);

-- layer0_node1_MUX[bit_math_h_l29_c3_432d]
signal layer0_node1_MUX_bit_math_h_l29_c3_432d_cond : unsigned(0 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue : unsigned(31 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse : unsigned(31 downto 0);
signal layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output : unsigned(31 downto 0);

-- layer0_node2_MUX[bit_math_h_l40_c3_775a]
signal layer0_node2_MUX_bit_math_h_l40_c3_775a_cond : unsigned(0 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue : unsigned(31 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse : unsigned(31 downto 0);
signal layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output : unsigned(31 downto 0);

-- layer0_node3_MUX[bit_math_h_l51_c3_00a7]
signal layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond : unsigned(0 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue : unsigned(31 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse : unsigned(31 downto 0);
signal layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output : unsigned(31 downto 0);

-- layer0_node4_MUX[bit_math_h_l62_c3_0480]
signal layer0_node4_MUX_bit_math_h_l62_c3_0480_cond : unsigned(0 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue : unsigned(31 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse : unsigned(31 downto 0);
signal layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output : unsigned(31 downto 0);

-- layer0_node5_MUX[bit_math_h_l73_c3_6955]
signal layer0_node5_MUX_bit_math_h_l73_c3_6955_cond : unsigned(0 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue : unsigned(31 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse : unsigned(31 downto 0);
signal layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output : unsigned(31 downto 0);

-- layer0_node6_MUX[bit_math_h_l84_c3_188d]
signal layer0_node6_MUX_bit_math_h_l84_c3_188d_cond : unsigned(0 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue : unsigned(31 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse : unsigned(31 downto 0);
signal layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output : unsigned(31 downto 0);

-- layer0_node7_MUX[bit_math_h_l95_c3_ee26]
signal layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond : unsigned(0 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue : unsigned(31 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse : unsigned(31 downto 0);
signal layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output : unsigned(31 downto 0);

-- layer1_node0_MUX[bit_math_h_l112_c3_e606]
signal layer1_node0_MUX_bit_math_h_l112_c3_e606_cond : unsigned(0 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue : unsigned(31 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse : unsigned(31 downto 0);
signal layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output : unsigned(31 downto 0);

-- layer1_node1_MUX[bit_math_h_l123_c3_af44]
signal layer1_node1_MUX_bit_math_h_l123_c3_af44_cond : unsigned(0 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue : unsigned(31 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse : unsigned(31 downto 0);
signal layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output : unsigned(31 downto 0);

-- layer1_node2_MUX[bit_math_h_l134_c3_d958]
signal layer1_node2_MUX_bit_math_h_l134_c3_d958_cond : unsigned(0 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue : unsigned(31 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse : unsigned(31 downto 0);
signal layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output : unsigned(31 downto 0);

-- layer1_node3_MUX[bit_math_h_l145_c3_6197]
signal layer1_node3_MUX_bit_math_h_l145_c3_6197_cond : unsigned(0 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue : unsigned(31 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse : unsigned(31 downto 0);
signal layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output : unsigned(31 downto 0);

-- layer2_node0_MUX[bit_math_h_l162_c3_9962]
signal layer2_node0_MUX_bit_math_h_l162_c3_9962_cond : unsigned(0 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue : unsigned(31 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse : unsigned(31 downto 0);
signal layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output : unsigned(31 downto 0);

-- layer2_node1_MUX[bit_math_h_l173_c3_92dc]
signal layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond : unsigned(0 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue : unsigned(31 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse : unsigned(31 downto 0);
signal layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output : unsigned(31 downto 0);

-- layer3_node0_MUX[bit_math_h_l190_c3_05a1]
signal layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond : unsigned(0 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue : unsigned(31 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse : unsigned(31 downto 0);
signal layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output : unsigned(31 downto 0);

function uint4_0_0( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(0- i);
      end loop;
return return_output;
end function;

function uint4_1_1( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(1- i);
      end loop;
return return_output;
end function;

function uint4_2_2( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(2- i);
      end loop;
return return_output;
end function;

function uint4_3_3( x : unsigned) return unsigned is
--variable x : unsigned(3 downto 0);
  variable return_output : unsigned(0 downto 0);
begin
for i in 0 to return_output'length-1 loop
        return_output(i) := x(3- i);
      end loop;
return return_output;
end function;


begin

-- SUBMODULE INSTANCES 
-- layer0_node0_MUX_bit_math_h_l18_c3_2607 : 0 clocks latency
layer0_node0_MUX_bit_math_h_l18_c3_2607 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node0_MUX_bit_math_h_l18_c3_2607_cond,
layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue,
layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse,
layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output);

-- layer0_node1_MUX_bit_math_h_l29_c3_432d : 0 clocks latency
layer0_node1_MUX_bit_math_h_l29_c3_432d : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node1_MUX_bit_math_h_l29_c3_432d_cond,
layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue,
layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse,
layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output);

-- layer0_node2_MUX_bit_math_h_l40_c3_775a : 0 clocks latency
layer0_node2_MUX_bit_math_h_l40_c3_775a : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node2_MUX_bit_math_h_l40_c3_775a_cond,
layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue,
layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse,
layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output);

-- layer0_node3_MUX_bit_math_h_l51_c3_00a7 : 0 clocks latency
layer0_node3_MUX_bit_math_h_l51_c3_00a7 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond,
layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue,
layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse,
layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output);

-- layer0_node4_MUX_bit_math_h_l62_c3_0480 : 0 clocks latency
layer0_node4_MUX_bit_math_h_l62_c3_0480 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node4_MUX_bit_math_h_l62_c3_0480_cond,
layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue,
layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse,
layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output);

-- layer0_node5_MUX_bit_math_h_l73_c3_6955 : 0 clocks latency
layer0_node5_MUX_bit_math_h_l73_c3_6955 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node5_MUX_bit_math_h_l73_c3_6955_cond,
layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue,
layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse,
layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output);

-- layer0_node6_MUX_bit_math_h_l84_c3_188d : 0 clocks latency
layer0_node6_MUX_bit_math_h_l84_c3_188d : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node6_MUX_bit_math_h_l84_c3_188d_cond,
layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue,
layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse,
layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output);

-- layer0_node7_MUX_bit_math_h_l95_c3_ee26 : 0 clocks latency
layer0_node7_MUX_bit_math_h_l95_c3_ee26 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond,
layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue,
layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse,
layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output);

-- layer1_node0_MUX_bit_math_h_l112_c3_e606 : 0 clocks latency
layer1_node0_MUX_bit_math_h_l112_c3_e606 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer1_node0_MUX_bit_math_h_l112_c3_e606_cond,
layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue,
layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse,
layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output);

-- layer1_node1_MUX_bit_math_h_l123_c3_af44 : 0 clocks latency
layer1_node1_MUX_bit_math_h_l123_c3_af44 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer1_node1_MUX_bit_math_h_l123_c3_af44_cond,
layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue,
layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse,
layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output);

-- layer1_node2_MUX_bit_math_h_l134_c3_d958 : 0 clocks latency
layer1_node2_MUX_bit_math_h_l134_c3_d958 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer1_node2_MUX_bit_math_h_l134_c3_d958_cond,
layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue,
layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse,
layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output);

-- layer1_node3_MUX_bit_math_h_l145_c3_6197 : 0 clocks latency
layer1_node3_MUX_bit_math_h_l145_c3_6197 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer1_node3_MUX_bit_math_h_l145_c3_6197_cond,
layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue,
layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse,
layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output);

-- layer2_node0_MUX_bit_math_h_l162_c3_9962 : 0 clocks latency
layer2_node0_MUX_bit_math_h_l162_c3_9962 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer2_node0_MUX_bit_math_h_l162_c3_9962_cond,
layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue,
layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse,
layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output);

-- layer2_node1_MUX_bit_math_h_l173_c3_92dc : 0 clocks latency
layer2_node1_MUX_bit_math_h_l173_c3_92dc : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond,
layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue,
layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse,
layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output);

-- layer3_node0_MUX_bit_math_h_l190_c3_05a1 : 0 clocks latency
layer3_node0_MUX_bit_math_h_l190_c3_05a1 : entity work.MUX_uint1_t_uint32_t_uint32_t_0CLK_de264c78 port map (
layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond,
layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue,
layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse,
layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 sel,
 in0,
 in1,
 in2,
 in3,
 in4,
 in5,
 in6,
 in7,
 in8,
 in9,
 in10,
 in11,
 in12,
 in13,
 in14,
 in15,
 -- All submodule outputs
 layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output,
 layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output,
 layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output,
 layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output,
 layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output,
 layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output,
 layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output,
 layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output,
 layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output,
 layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output,
 layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output,
 layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output,
 layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output,
 layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output,
 layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : unsigned(31 downto 0);
 variable VAR_sel : unsigned(3 downto 0);
 variable VAR_in0 : unsigned(31 downto 0);
 variable VAR_in1 : unsigned(31 downto 0);
 variable VAR_in2 : unsigned(31 downto 0);
 variable VAR_in3 : unsigned(31 downto 0);
 variable VAR_in4 : unsigned(31 downto 0);
 variable VAR_in5 : unsigned(31 downto 0);
 variable VAR_in6 : unsigned(31 downto 0);
 variable VAR_in7 : unsigned(31 downto 0);
 variable VAR_in8 : unsigned(31 downto 0);
 variable VAR_in9 : unsigned(31 downto 0);
 variable VAR_in10 : unsigned(31 downto 0);
 variable VAR_in11 : unsigned(31 downto 0);
 variable VAR_in12 : unsigned(31 downto 0);
 variable VAR_in13 : unsigned(31 downto 0);
 variable VAR_in14 : unsigned(31 downto 0);
 variable VAR_in15 : unsigned(31 downto 0);
 variable VAR_sel0 : unsigned(0 downto 0);
 variable VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output : unsigned(0 downto 0);
 variable VAR_layer0_node0 : unsigned(31 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_cond : unsigned(0 downto 0);
 variable VAR_layer0_node1 : unsigned(31 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node2 : unsigned(31 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_cond : unsigned(0 downto 0);
 variable VAR_layer0_node3 : unsigned(31 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond : unsigned(0 downto 0);
 variable VAR_layer0_node4 : unsigned(31 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_cond : unsigned(0 downto 0);
 variable VAR_layer0_node5 : unsigned(31 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_cond : unsigned(0 downto 0);
 variable VAR_layer0_node6 : unsigned(31 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_cond : unsigned(0 downto 0);
 variable VAR_layer0_node7 : unsigned(31 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue : unsigned(31 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse : unsigned(31 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output : unsigned(31 downto 0);
 variable VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond : unsigned(0 downto 0);
 variable VAR_sel1 : unsigned(0 downto 0);
 variable VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output : unsigned(0 downto 0);
 variable VAR_layer1_node0 : unsigned(31 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue : unsigned(31 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse : unsigned(31 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output : unsigned(31 downto 0);
 variable VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_cond : unsigned(0 downto 0);
 variable VAR_layer1_node1 : unsigned(31 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue : unsigned(31 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse : unsigned(31 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output : unsigned(31 downto 0);
 variable VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_cond : unsigned(0 downto 0);
 variable VAR_layer1_node2 : unsigned(31 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue : unsigned(31 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse : unsigned(31 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output : unsigned(31 downto 0);
 variable VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_cond : unsigned(0 downto 0);
 variable VAR_layer1_node3 : unsigned(31 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue : unsigned(31 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse : unsigned(31 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output : unsigned(31 downto 0);
 variable VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_cond : unsigned(0 downto 0);
 variable VAR_sel2 : unsigned(0 downto 0);
 variable VAR_uint4_2_2_bit_math_h_l158_c10_cac1_return_output : unsigned(0 downto 0);
 variable VAR_layer2_node0 : unsigned(31 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue : unsigned(31 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse : unsigned(31 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output : unsigned(31 downto 0);
 variable VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_cond : unsigned(0 downto 0);
 variable VAR_layer2_node1 : unsigned(31 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue : unsigned(31 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse : unsigned(31 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output : unsigned(31 downto 0);
 variable VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond : unsigned(0 downto 0);
 variable VAR_sel3 : unsigned(0 downto 0);
 variable VAR_uint4_3_3_bit_math_h_l186_c10_c591_return_output : unsigned(0 downto 0);
 variable VAR_layer3_node0 : unsigned(31 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue : unsigned(31 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse : unsigned(31 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output : unsigned(31 downto 0);
 variable VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond : unsigned(0 downto 0);
begin

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_sel := sel;
     VAR_in0 := in0;
     VAR_in1 := in1;
     VAR_in2 := in2;
     VAR_in3 := in3;
     VAR_in4 := in4;
     VAR_in5 := in5;
     VAR_in6 := in6;
     VAR_in7 := in7;
     VAR_in8 := in8;
     VAR_in9 := in9;
     VAR_in10 := in10;
     VAR_in11 := in11;
     VAR_in12 := in12;
     VAR_in13 := in13;
     VAR_in14 := in14;
     VAR_in15 := in15;

     -- Submodule level 0
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse := VAR_in0;
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue := VAR_in1;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse := VAR_in10;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue := VAR_in11;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse := VAR_in12;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue := VAR_in13;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse := VAR_in14;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue := VAR_in15;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse := VAR_in2;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue := VAR_in3;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse := VAR_in4;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue := VAR_in5;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse := VAR_in6;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue := VAR_in7;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse := VAR_in8;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue := VAR_in9;
     -- uint4_3_3[bit_math_h_l186_c10_c591] LATENCY=0
     VAR_uint4_3_3_bit_math_h_l186_c10_c591_return_output := uint4_3_3(
     VAR_sel);

     -- uint4_0_0[bit_math_h_l14_c10_6f73] LATENCY=0
     VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output := uint4_0_0(
     VAR_sel);

     -- uint4_2_2[bit_math_h_l158_c10_cac1] LATENCY=0
     VAR_uint4_2_2_bit_math_h_l158_c10_cac1_return_output := uint4_2_2(
     VAR_sel);

     -- uint4_1_1[bit_math_h_l108_c10_b4e9] LATENCY=0
     VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output := uint4_1_1(
     VAR_sel);

     -- Submodule level 1
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond := VAR_uint4_0_0_bit_math_h_l14_c10_6f73_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_cond := VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_cond := VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_cond := VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_cond := VAR_uint4_1_1_bit_math_h_l108_c10_b4e9_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_cond := VAR_uint4_2_2_bit_math_h_l158_c10_cac1_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond := VAR_uint4_2_2_bit_math_h_l158_c10_cac1_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond := VAR_uint4_3_3_bit_math_h_l186_c10_c591_return_output;
     -- layer0_node5_MUX[bit_math_h_l73_c3_6955] LATENCY=0
     -- Inputs
     layer0_node5_MUX_bit_math_h_l73_c3_6955_cond <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_cond;
     layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iftrue;
     layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse <= VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_iffalse;
     -- Outputs
     VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output := layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output;

     -- layer0_node1_MUX[bit_math_h_l29_c3_432d] LATENCY=0
     -- Inputs
     layer0_node1_MUX_bit_math_h_l29_c3_432d_cond <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_cond;
     layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iftrue;
     layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse <= VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_iffalse;
     -- Outputs
     VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output := layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output;

     -- layer0_node4_MUX[bit_math_h_l62_c3_0480] LATENCY=0
     -- Inputs
     layer0_node4_MUX_bit_math_h_l62_c3_0480_cond <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_cond;
     layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iftrue;
     layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse <= VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_iffalse;
     -- Outputs
     VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output := layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output;

     -- layer0_node3_MUX[bit_math_h_l51_c3_00a7] LATENCY=0
     -- Inputs
     layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_cond;
     layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iftrue;
     layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse <= VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_iffalse;
     -- Outputs
     VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output := layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output;

     -- layer0_node6_MUX[bit_math_h_l84_c3_188d] LATENCY=0
     -- Inputs
     layer0_node6_MUX_bit_math_h_l84_c3_188d_cond <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_cond;
     layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iftrue;
     layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse <= VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_iffalse;
     -- Outputs
     VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output := layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output;

     -- layer0_node2_MUX[bit_math_h_l40_c3_775a] LATENCY=0
     -- Inputs
     layer0_node2_MUX_bit_math_h_l40_c3_775a_cond <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_cond;
     layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iftrue;
     layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse <= VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_iffalse;
     -- Outputs
     VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output := layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output;

     -- layer0_node0_MUX[bit_math_h_l18_c3_2607] LATENCY=0
     -- Inputs
     layer0_node0_MUX_bit_math_h_l18_c3_2607_cond <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_cond;
     layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iftrue;
     layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse <= VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_iffalse;
     -- Outputs
     VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output := layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output;

     -- layer0_node7_MUX[bit_math_h_l95_c3_ee26] LATENCY=0
     -- Inputs
     layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_cond;
     layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iftrue;
     layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse <= VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_iffalse;
     -- Outputs
     VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output := layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output;

     -- Submodule level 2
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse := VAR_layer0_node0_MUX_bit_math_h_l18_c3_2607_return_output;
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue := VAR_layer0_node1_MUX_bit_math_h_l29_c3_432d_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse := VAR_layer0_node2_MUX_bit_math_h_l40_c3_775a_return_output;
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue := VAR_layer0_node3_MUX_bit_math_h_l51_c3_00a7_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse := VAR_layer0_node4_MUX_bit_math_h_l62_c3_0480_return_output;
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue := VAR_layer0_node5_MUX_bit_math_h_l73_c3_6955_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse := VAR_layer0_node6_MUX_bit_math_h_l84_c3_188d_return_output;
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue := VAR_layer0_node7_MUX_bit_math_h_l95_c3_ee26_return_output;
     -- layer1_node1_MUX[bit_math_h_l123_c3_af44] LATENCY=0
     -- Inputs
     layer1_node1_MUX_bit_math_h_l123_c3_af44_cond <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_cond;
     layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iftrue;
     layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse <= VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_iffalse;
     -- Outputs
     VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output := layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output;

     -- layer1_node3_MUX[bit_math_h_l145_c3_6197] LATENCY=0
     -- Inputs
     layer1_node3_MUX_bit_math_h_l145_c3_6197_cond <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_cond;
     layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iftrue;
     layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse <= VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_iffalse;
     -- Outputs
     VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output := layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output;

     -- layer1_node0_MUX[bit_math_h_l112_c3_e606] LATENCY=0
     -- Inputs
     layer1_node0_MUX_bit_math_h_l112_c3_e606_cond <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_cond;
     layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iftrue;
     layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse <= VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_iffalse;
     -- Outputs
     VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output := layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output;

     -- layer1_node2_MUX[bit_math_h_l134_c3_d958] LATENCY=0
     -- Inputs
     layer1_node2_MUX_bit_math_h_l134_c3_d958_cond <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_cond;
     layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iftrue;
     layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse <= VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_iffalse;
     -- Outputs
     VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output := layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output;

     -- Submodule level 3
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse := VAR_layer1_node0_MUX_bit_math_h_l112_c3_e606_return_output;
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue := VAR_layer1_node1_MUX_bit_math_h_l123_c3_af44_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse := VAR_layer1_node2_MUX_bit_math_h_l134_c3_d958_return_output;
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue := VAR_layer1_node3_MUX_bit_math_h_l145_c3_6197_return_output;
     -- layer2_node1_MUX[bit_math_h_l173_c3_92dc] LATENCY=0
     -- Inputs
     layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_cond;
     layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iftrue;
     layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse <= VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_iffalse;
     -- Outputs
     VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output := layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output;

     -- layer2_node0_MUX[bit_math_h_l162_c3_9962] LATENCY=0
     -- Inputs
     layer2_node0_MUX_bit_math_h_l162_c3_9962_cond <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_cond;
     layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iftrue;
     layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse <= VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_iffalse;
     -- Outputs
     VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output := layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output;

     -- Submodule level 4
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse := VAR_layer2_node0_MUX_bit_math_h_l162_c3_9962_return_output;
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue := VAR_layer2_node1_MUX_bit_math_h_l173_c3_92dc_return_output;
     -- layer3_node0_MUX[bit_math_h_l190_c3_05a1] LATENCY=0
     -- Inputs
     layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_cond;
     layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iftrue;
     layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse <= VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_iffalse;
     -- Outputs
     VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output := layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output;

     -- Submodule level 5
     VAR_return_output := VAR_layer3_node0_MUX_bit_math_h_l190_c3_05a1_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
