-- Timing params:
--   Fixed?: False
--   Pipeline Slices: []
--   Input regs?: False
--   Output regs?: False
library std;
use std.textio.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.float_pkg.all;
use work.c_structs_pkg.all;
-- Submodules: 17
entity work_0CLK_83e31706 is
port(
 inputs : in work_inputs_t;
 return_output : out work_outputs_t);
end work_0CLK_83e31706;
architecture arch of work_0CLK_83e31706 is
-- Types and such
-- Declarations
attribute mark_debug : string;
constant ADDED_PIPELINE_LATENCY : integer := 0;
-- All of the wires/regs in function
-- Each function instance gets signals
-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_4439]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_345f]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_b777]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_63a6]
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_0ea4]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_439b]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_f436]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output : signed(16 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_4806]
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left : signed(7 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right : signed(15 downto 0);
signal FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output : signed(16 downto 0);

function CONST_REF_RD_work_outputs_t_work_outputs_t_c871( ref_toks_0 : signed;
 ref_toks_1 : signed;
 ref_toks_2 : signed;
 ref_toks_3 : signed) return work_outputs_t is
 
  variable base : work_outputs_t; 
  variable return_output : work_outputs_t;
begin
      base.result(0)(0) := ref_toks_0;
      base.result(0)(1) := ref_toks_1;
      base.result(1)(0) := ref_toks_2;
      base.result(1)(1) := ref_toks_3;

      return_output := base;
      return return_output; 
end function;


begin

-- SUBMODULE INSTANCES 
-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right,
FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9 : entity work.BIN_OP_INFERRED_MULT_int8_t_int8_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output);

-- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806 : 0 clocks latency
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806 : entity work.BIN_OP_PLUS_int8_t_int16_t_0CLK_de264c78 port map (
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right,
FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output);



-- Combinatorial process for pipeline stages
process (
 -- Inputs
 inputs,
 -- All submodule outputs
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output,
 FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output)
is 
 -- All of the wires in function
 variable VAR_CLOCK_ENABLE : unsigned(0 downto 0);
 variable VAR_return_output : work_outputs_t;
 variable VAR_inputs : work_inputs_t;
 variable VAR_outputs : work_outputs_t;
 variable VAR_i : unsigned(31 downto 0);
 variable VAR_j : unsigned(31 downto 0);
 variable VAR_k : unsigned(31 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_0_0_work_h_l67_c13_2db5 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_0_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_0_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_0_1_work_h_l67_c13_2db5 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_1_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_1_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_1_0_work_h_l67_c13_2db5 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_0_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_0_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_1_1_work_h_l67_c13_2db5 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_1_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output : signed(16 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_1_work_h_l70_c17_f9b8 : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right : signed(7 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right : signed(15 downto 0);
 variable VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output : signed(16 downto 0);
 variable VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_adba_return_output : work_outputs_t;
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_578c_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_6755_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_f1dc_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_9a22_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_4d72_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_bdea_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_f67e_return_output : signed(7 downto 0);
 variable VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_290c_return_output : signed(7 downto 0);
begin
 -- Constants and things derived from constants alone
     -- Submodule level 0
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_1_1_work_h_l67_c13_2db5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_1_1_work_h_l67_c13_2db5;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_0_1_work_h_l67_c13_2db5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_outputs_result_0_1_work_h_l67_c13_2db5;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_1_0_work_h_l67_c13_2db5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_1_0_work_h_l67_c13_2db5;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_0_0_work_h_l67_c13_2db5 := signed(std_logic_vector(resize(to_unsigned(0, 1), 8)));
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_outputs_result_0_0_work_h_l67_c13_2db5;

 -- Loop to construct simultaneous register transfers for each of the pipeline stages
 -- LATENCY=0 is combinational Logic
 for STAGE in 0 to ADDED_PIPELINE_LATENCY loop
   if STAGE = 0 then
     -- Mux in inputs
     VAR_inputs := inputs;

     -- Submodule level 0
     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d[work_h_l70_c41_e4cb]_DUPLICATE_f1dc LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_f1dc_return_output := VAR_inputs.matrix0(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d[work_h_l70_c41_e4cb]_DUPLICATE_290c LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_290c_return_output := VAR_inputs.matrix0(1)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d[work_h_l70_c64_a8ec]_DUPLICATE_9a22 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_9a22_return_output := VAR_inputs.matrix1(1)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d[work_h_l70_c64_a8ec]_DUPLICATE_6755 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_6755_return_output := VAR_inputs.matrix1(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d[work_h_l70_c41_e4cb]_DUPLICATE_578c LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_578c_return_output := VAR_inputs.matrix0(0)(0);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d[work_h_l70_c64_a8ec]_DUPLICATE_bdea LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_bdea_return_output := VAR_inputs.matrix1(1)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d[work_h_l70_c64_a8ec]_DUPLICATE_4d72 LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_4d72_return_output := VAR_inputs.matrix1(0)(1);

     -- CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d[work_h_l70_c41_e4cb]_DUPLICATE_f67e LATENCY=0
     VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_f67e_return_output := VAR_inputs.matrix0(1)(0);

     -- Submodule level 1
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_578c_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_578c_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_f1dc_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_0_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_f1dc_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_f67e_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_0_d41d_work_h_l70_c41_e4cb_DUPLICATE_f67e_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_290c_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix0_1_1_d41d_work_h_l70_c41_e4cb_DUPLICATE_290c_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_6755_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_6755_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_4d72_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_0_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_4d72_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_9a22_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_0_d41d_work_h_l70_c64_a8ec_DUPLICATE_9a22_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_bdea_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right := VAR_CONST_REF_RD_int8_t_work_inputs_t_matrix1_1_1_d41d_work_h_l70_c64_a8ec_DUPLICATE_bdea_return_output;
     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT[work_h_l70_c41_27c9] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;

     -- Submodule level 2
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_INFERRED_MULT_work_h_l70_c41_27c9_return_output;
     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_4439] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_b777] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_f436] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS[work_h_l70_c17_0ea4] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output;

     -- Submodule level 3
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_0_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_4439_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_1_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_b777_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_0_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_0ea4_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_1_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_BIN_OP_PLUS_work_h_l70_c17_f436_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_0_work_h_l70_c17_f9b8;
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left := VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_0_1_work_h_l70_c17_f9b8;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_0_work_h_l70_c17_f9b8;
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left := VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_0_outputs_result_1_1_work_h_l70_c17_f9b8;
     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_4806] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_63a6] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_345f] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_left;
     FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output := FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output;

     -- FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS[work_h_l70_c17_439b] LATENCY=0
     -- Inputs
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_left;
     FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right <= VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_right;
     -- Outputs
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output := FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output;

     -- Submodule level 4
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_0_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_345f_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_1_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_63a6_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_0_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_439b_return_output, 8);
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_1_work_h_l70_c17_f9b8 := resize(VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_BIN_OP_PLUS_work_h_l70_c17_4806_return_output, 8);
     -- CONST_REF_RD_work_outputs_t_work_outputs_t_c871[work_h_l74_c12_adba] LATENCY=0
     VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_adba_return_output := CONST_REF_RD_work_outputs_t_work_outputs_t_c871(
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_0_work_h_l70_c17_f9b8,
     VAR_FOR_work_h_l63_c5_66c5_ITER_0_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_0_1_work_h_l70_c17_f9b8,
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_0_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_0_work_h_l70_c17_f9b8,
     VAR_FOR_work_h_l63_c5_66c5_ITER_1_FOR_work_h_l65_c9_063c_ITER_1_FOR_work_h_l68_c13_6aa1_ITER_1_outputs_result_1_1_work_h_l70_c17_f9b8);

     -- Submodule level 5
     VAR_return_output := VAR_CONST_REF_RD_work_outputs_t_work_outputs_t_c871_work_h_l74_c12_adba_return_output;
     -- Last stage of pipeline return wire to return port/reg
     return_output <= VAR_return_output;
   end if;
 end loop;

end process;

end arch;
